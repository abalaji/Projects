library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.user_pkg.all;

entity dual_flop_h101 is
  port(
    clk1 : in  std_logic;
    clk2 : in  std_logic;
    rst  : in  std_logic;
    addr : in  std_logic_vector(31 downto 0);
    en   : in  std_logic;
    wen  : in  std_logic;
    din  : in  std_logic_vector(31 downto 0);
    dout : out std_logic_vector(31 downto 0)
    );

  attribute dtinfo         : string;
  attribute dtinfo of clk1 : signal is "clk1";
  attribute dtinfo of clk2 : signal is "clk2";
  attribute dtinfo of rst  : signal  is "reset";
  attribute dtinfo of addr : signal is "usergroup, memmap";
end dual_flop_h101;

architecture STR of dual_flop_h101 is

  signal iterations         : std_logic_vector(31 downto 0);
  signal count              : std_logic_vector(31 downto 0);
  signal pulse              : std_logic;
  signal go                 : std_logic;
  signal done, done_delayed : std_logic;
  signal dest_rst           : std_logic;
  signal ff1_out, ff2_out, dfs_out : std_logic;
begin

  -----------------------------------------------------------------------------
  -- Clock domain 1

  U_GLUE_LOGIC : entity work.glue_logic
    port map (
      clk        => clk1,
      rst        => rst,
      addr       => addr,
      en         => en,
      wen        => wen,
      din        => din,
      dout       => dout,
      go         => go,
      iterations => iterations,
      count      => count,
      done       => done_delayed);

  -- source generates "iterations" numbers of pulses  
  U_SOURCE : entity work.source
    generic map (
      clk_in_freq      => C_SRC_DEST_CLK_RATIO,
      clk_out_freq     => 1,
      iterations_width => 32)
    port map (
      clk              => clk1,
      rst              => rst,
      iterations       => iterations,
      go               => go,
      done             => done,
      output           => pulse);

  -- this delays the done signal to make sure that the destination domain has
  -- time to see the final pulse
  U_DELAY : entity work.delay
    generic map (
      cycles    => 10,                  -- assume 10 cycles is plenty for sync
      width     => 1)
    port map (
      clk       => clk1,
      rst       => dest_rst,
      en        => C_1,
      input(0)  => done,
      output(0) => done_delayed);

  -----------------------------------------------------------------------------
  -- Clock domain 2

  -- Dest is a counter in the destination clock domain that counts the number
  -- of times that the input signal transitions from 0 to 1. The input signal
  -- is generated by the pulses in the source domain.

  U_DEST : entity work.dest
    generic map (
      width  => 32)
    port map (
      clk    => clk2,
      rst    => dest_rst,
		input => dfs_out,
      --input  => pulse,                  -- INCORRECT: not synchronized, will go metastable
      output => count);

  -- simple way to make sure dest counter is cleared every time
  dest_rst <= go or rst;

  -----------------------------------------------------------------------------
  -- CDC

  -- TODO: Instantiate a dual flop synchronizer to properly synchronize the
  -- pulse signal that crosses domain 1 to domain 2. You will also need to make
  -- minor corrections to the other parts of the code.

	U_FF1 : entity work.reg
	generic map (
				width => 1)
			port map ( clk => clk1,
						rst => rst,
						en => C_1,
						input(0) => pulse,
						output(0) => ff1_out);

	U_FF2 : entity work.reg
	generic map(
				width => 1)
			port map ( clk => clk2,
						rst => dest_rst,
						en => C_1,
						input(0) => ff1_out,
						output(0) => ff2_out);
						
	U_FF3 : entity work.reg
	generic map(
				width => 1)
			port map ( clk => clk2,
						rst => dest_rst,
						en => C_1,
						input(0) => ff2_out,
						output(0) => dfs_out);
						
  -- There is actually another synchronization problem with this code that
  -- you are not required to fix in this part. However, you should try to
  -- identify it.

end STR;
