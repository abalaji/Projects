-- Greg Stitt
-- University of Florida
-- EEL 5934/4930 Reconfigurable Computing
--
-- File: ctrl.vhd
--
-- Description: This file implements the controller for the Fibonacci
-- calculator
--
-- Comments: The FSM was kept simple for ease of understanding. It can
-- certainly be optimized if you want to put in the extra effort.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ctrl is
  port( clk, rst, go : in  std_logic;
        done         : out std_logic;

        -- control signals used/generated by the datapath
        i_sel, x_sel, y_sel               : out std_logic;
        i_ld, x_ld, y_ld, n_ld, result_ld : out std_logic;
        i_le_n                            : in  std_logic );
end ctrl;

architecture bhv of ctrl is

  type STATE_TYPE is (START, WAIT_0, WAIT_1, INIT, LOOP_COND,
                      LOOP_BODY, RESULT);
  signal state, next_state   : STATE_TYPE;
  signal done_s, next_done_s : std_logic;

begin

  -- state register
  process (clk, rst)
  begin
    if (rst = '1') then
      state  <= START;
      done_s <= '0';
    elsif (clk = '1' and clk'event) then
      state  <= next_state;
      done_s <= next_done_s;
    end if;
  end process;

  -- next state logic
  process( go, i_le_n, state, done_s )
  begin

    i_sel <= '-';
    x_sel <= '-';
    y_sel <= '-';
    i_ld  <= '-';
    x_ld  <= '-';
    y_ld  <= '-';
    n_ld  <= '-';
    result_ld <= '-';
    
    next_done_s <= done_s;
    next_state  <= state;

    case state is
      when START =>

        result_ld <= '0';

        if (go = '0') then
          next_state <= WAIT_1;
        end if;

      when WAIT_1 =>

        result_ld <= '0';

        if (go = '1') then
          next_done_s <= '0';
          next_state  <= INIT;
        end if;

      when INIT =>

        i_sel     <= '1';
        x_sel     <= '1';
        y_sel     <= '1';
        i_ld      <= '1';
        x_ld      <= '1';
        y_ld      <= '1';
        n_ld      <= '1';
        result_ld <= '0';

        next_state <= LOOP_COND;

      when LOOP_COND =>

        i_ld      <= '0';
        x_ld      <= '0';
        y_ld      <= '0';
        n_ld      <= '0';
        result_ld <= '0';

        if (i_le_n = '1') then
          next_state <= LOOP_BODY;
        else
          next_state <= RESULT;
        end if;

      when LOOP_BODY =>

        i_sel     <= '0';
        x_sel     <= '0';
        y_sel     <= '0';
        i_ld      <= '1';
        x_ld      <= '1';
        y_ld      <= '1';
        n_ld      <= '0';
        result_ld <= '0';

        next_state <= LOOP_COND;

      when RESULT =>
        next_done_s  <= '1';
        result_ld  <= '1';
        next_state <= WAIT_0;

      when WAIT_0 =>

        result_ld <= '0';

        if (go = '0') then
          next_state <= WAIT_1;
        end if;

      when others => null;
    end case;
  end process;

  done <= done_s;
  
end bhv;
